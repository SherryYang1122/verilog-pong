`timescale 1ns / 1ps
module vsync_unit(
    );


endmodule

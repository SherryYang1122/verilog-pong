`timescale 1ns / 1ps
module graph_unit(
    );


endmodule
